library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testbench_up_down_counter is
end entity;

architecture is
	signal 
