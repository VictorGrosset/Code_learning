library IEEE;
use IEEE.std_logic_1164.all;



entity testbench_deco7seg is
end entity;



architecture ar of testbench_deco7seg is


begin



end architecture;
